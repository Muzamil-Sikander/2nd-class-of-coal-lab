//  Combinational Circuit
module C_Circuit (a,b,c,o);

//  declaring inputs and output
 input a;
 input b;
 input c;

 output o;

//  Interm Wire

wire X ;

assign x = a | b ;
assign o = x & c ;






endmodule

